module x87_format; endmodule
