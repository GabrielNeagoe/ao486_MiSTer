module x87_format(input wire clk,input wire rst); endmodule
