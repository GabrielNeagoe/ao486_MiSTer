module x87_divsqrt(input wire clk,input wire rst); endmodule
